/////////////////////////////////////////////////////////////////////
// Design unit: rotation_cordic
//            :
// File name  : rotation_cordic.sv
//            :
//            :
// Replace <ecsid> with your ECS ID below
//
// Author     : <ecsid>@ecs.soton.ac.uk
/////////////////////////////////////////////////////////////////////

// Do not change this next line

module rotation_cordic(output logic data_out_rot, output logic [15:0] xprime, output logic [15:0] yprime, input logic [15:0] x,input logic [15:0] y,input logic [15:0] theta,input logic Clk, Reset, Start);


// Include your design here

endmodule
