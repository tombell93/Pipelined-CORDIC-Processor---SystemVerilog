/////////////////////////////////////////////////////////////////////
// Design unit: cordic
//            :
// File name  : cordic_top.sv
//            :
//            :
// Replace <ecsid> with your ECS ID below
//
// Author     : <ecsid>@ecs.soton.ac.uk
/////////////////////////////////////////////////////////////////////

// Do not change this next line

module cordic_top (output logic data_out, output logic [15:0] X, output logic [15:0] Y, 
input logic [15:0] x, input logic [15:0] y, input logic [15:0] a, input logic [15:0] b,input logic Clk, Reset, Start);

// Include your top level architecture here

endmodule


