/////////////////////////////////////////////////////////////////////
// Design unit: vector_cordic
//            :
// File name  : vector_cordic.sv
//            :
//            :
// Replace <ecsid> with your ECS ID below
//
// Author     : <ecsid>@ecs.soton.ac.uk
/////////////////////////////////////////////////////////////////////

// Do not change this next line

module vector_cordic(output logic data_out_vec, output logic [15:0] rootxy, output logic [15:0] atanba, input logic [15:0] x,input logic [15:0] y,input logic [15:0] z,input logic Clk, Reset, Start);


// Include your design here

endmodule

