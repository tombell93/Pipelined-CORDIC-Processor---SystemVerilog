library verilog;
use verilog.vl_types.all;
entity cordic_test is
    generic(
        CLK12_SPEED     : real    := 40.700000
    );
end cordic_test;
