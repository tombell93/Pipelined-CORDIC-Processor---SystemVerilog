library verilog;
use verilog.vl_types.all;
entity MODEL is
end MODEL;
